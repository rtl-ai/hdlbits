//15_vector3.v

module top_module (
    input  [4:0] a,
    b,
    c,
    d,
    e,
    f,
    output [7:0] w,
    x,
    y,
    z
);

  wire [31:0] w_concat;

  assign w_concat = {a[4:0], b[4:0], c[4:0], d[4:0], e[4:0], f[4:0], 2'b11};

  assign w = w_concat[31:24];
  assign x = w_concat[23:16];
  assign y = w_concat[15:8];
  assign z = w_concat[7:0];

endmodule
